module Set_Number_Controler  (
                                input wire clk,
                                input wire rst,
                                input wire buttonUp,
                                input wire buttonCentre,
                                input wire buttonDown,
                                input wire buttonLeft,
                                input wire buttonRight,
                                output reg up,
                                output reg set,
                                output reg down,
                                output reg left,
                                output reg right
                             );

  wire [1:0]    upEdge,
                centreEdge,
                downEdge,
                leftEdge,
                rightEdge;

  EdgeDetector upEdgeDetector(.clk(clk), .rst(rst), .signal(buttonUp), .detected(upEdge));
  EdgeDetector centreEdgeDetector(.clk(clk), .rst(rst), .signal(buttonCentre), .detected(centreEdge));
  EdgeDetector downEdgeDetector(.clk(clk), .rst(rst), .signal(buttonDown), .detected(downEdge));
  EdgeDetector leftEdgeDetector(.clk(clk), .rst(rst), .signal(buttonLeft), .detected(leftEdge));
  EdgeDetector rightEdgeDetector(.clk(clk), .rst(rst), .signal(buttonRight), .detected(rightEdge));
  
  always @(posedge clk, posedge rst) begin
    if (rst) begin
        up <= 0;
        down <= 0;
        left <= 0;
        right <= 0;
        
        set <= set;
    end
    else begin
        up <= (upEdge == 2'b01)? 1:0;
        down <= (downEdge == 2'b01)? 1:0;
        left <= (leftEdge == 2'b01)? 1:0;
        right <= (rightEdge == 2'b01)? 1:0;
        
        set <= (centreEdge == 2'b01)? ~set:set;
    end
  end

endmodule
